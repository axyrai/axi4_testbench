package axi_sequence_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
endpackage  
