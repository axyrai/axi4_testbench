package axi_master_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "../../globals/axi_globals_pkg.sv"
import axi_globals_pkg::*;
endpackage
