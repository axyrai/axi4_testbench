package axi_master_pkg;
 `include "uvm_macros.svh"
 import uvm_pkg::*;
 import axi_env_pkg::*;
 import axi_master_pkg::*;
 import axi_sequence_pkg::*;
endpackage
