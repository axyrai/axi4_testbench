package axi_env_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import axi_globals_pkg::*;
  import axi_master_pkg::*;

  `include "axi_master_environment.sv"
  `include "axi_master_scoreboard.sv"
endpackage
