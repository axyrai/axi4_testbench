package axi_env_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;

endpackage
