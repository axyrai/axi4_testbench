package axi_env_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
    `include "../master/axi_master_transaction.sv"
`include "axi_master_scoreboard.sv"
`include "../master/axi_master_agent.sv"

endpackage
