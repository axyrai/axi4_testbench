package axi_master_pkg;
  `include "uvm_macros.svh"
  `include "../../globals/axi_globals_pkg.sv"
  import uvm_pkg::*;
  import axi_globals_pkg::*;
endpackage
