package axi_master_pkg;
 `include "uvm_macros.svh"
 import uvm_pkg::*;
endpackage
